module ex16 (
    
);
// this module can support both signed extend and unsigned extend

endmodule //ex16