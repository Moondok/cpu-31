module decoder(
    input[4:0] waddr,
    output reg [31:0] one_hot_waddr
    );
    always @(*)
    begin
        begin
            case (waddr)
                5'b00000: one_hot_waddr=32'b00000000_00000000_00000000_00000001;
                5'b00001: one_hot_waddr=32'b00000000_00000000_00000000_00000010;
                5'b00010: one_hot_waddr=32'b00000000_00000000_00000000_00000100;
                5'b00011: one_hot_waddr=32'b00000000_00000000_00000000_00001000;
                5'b00100: one_hot_waddr=32'b00000000_00000000_00000000_00010000;
                5'b00100: one_hot_waddr=32'b00000000_00000000_00000000_00100000;
                5'b00110: one_hot_waddr=32'b00000000_00000000_00000000_01000000;
                5'b00111: one_hot_waddr=32'b00000000_00000000_00000000_10000000;
                5'b01000: one_hot_waddr=32'b00000000_00000000_00000001_00000000;
                5'b01001: one_hot_waddr=32'b00000000_00000000_00000010_00000000;
                5'b01010: one_hot_waddr=32'b00000000_00000000_00000100_00000000;
                5'b01011: one_hot_waddr=32'b00000000_00000000_00001000_00000000;
                5'b01100: one_hot_waddr=32'b00000000_00000000_00010000_00000000;
                5'b01101: one_hot_waddr=32'b00000000_00000000_00100000_00000000;
                5'b01110: one_hot_waddr=32'b00000000_00000000_01000000_00000000;
                5'b01111: one_hot_waddr=32'b00000000_00000000_10000000_00000000;
                5'b10000: one_hot_waddr=32'b00000000_00000001_00000000_00000000;
                5'b10001: one_hot_waddr=32'b00000000_00000010_00000000_00000000;
                5'b10010: one_hot_waddr=32'b00000000_00000100_00000000_00000000;
                5'b10011: one_hot_waddr=32'b00000000_00001000_00000000_00000000;
                5'b10100: one_hot_waddr=32'b00000000_00010000_00000000_00000000;
                5'b10101: one_hot_waddr=32'b00000000_00100000_00000000_00000000;
                5'b10110: one_hot_waddr=32'b00000000_01000000_00000000_00000000;
                5'b10111: one_hot_waddr=32'b00000000_10000000_00000000_00000000;
                5'b11000: one_hot_waddr=32'b00000001_00000000_00000000_00000000;
                5'b11001: one_hot_waddr=32'b00000010_00000000_00000000_00000000;
                5'b11010: one_hot_waddr=32'b00000100_00000000_00000000_00000000;
                5'b11011: one_hot_waddr=32'b00001000_00000000_00000000_00000000;
                5'b11100: one_hot_waddr=32'b00010000_00000000_00000000_00000000;
                5'b11101: one_hot_waddr=32'b00100000_00000000_00000000_00000000;
                5'b11110: one_hot_waddr=32'b01000000_00000000_00000000_00000000;
                5'b11111: one_hot_waddr=32'b10000000_00000000_00000000_00000000;
                //5'b00010: one_hot_waddr=32'b00000000_00000000_00000000_00000010;
                
            endcase
        end
    end
endmodule