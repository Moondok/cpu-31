module controller (
    input [31:0] decoded_instr,
    output dmem_r,
    output dmem_w,
    output regfile_w,
    output [3:0] alu_control
);

endmodule //controller