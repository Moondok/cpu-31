module instrument_decoder (
    input [31:0] raw_instruction,
    output reg[31:0] code
);
// here we translate mips 32 instrument to one hot code
wire [11:0] tmp={raw_instruction[31:26],raw_instruction[5:0]};

// we transform mips instruction into one-hot code to generate control signal
always @(*) 
begin
    casex (tmp)
    //R-type
        12'b000000_100000: code<=32'b00000000_00000000_00000000_00000001;
        12'b000000_100001: code<=32'b00000000_00000000_00000000_00000010;
        12'b000000_100010: code<=32'b00000000_00000000_00000000_00000100;
        12'b000000_100011: code<=32'b00000000_00000000_00000000_00001000;
        12'b000000_100100: code<=32'b00000000_00000000_00000000_00010000;
        12'b000000_100101: code<=32'b00000000_00000000_00000000_00100000;
        12'b000000_100110: code<=32'b00000000_00000000_00000000_01000000;
        12'b000000_100111: code<=32'b00000000_00000000_00000000_10000000;
        12'b000000_101010: code<=32'b00000000_00000000_00000001_00000000;
        12'b000000_101011: code<=32'b00000000_00000000_00000010_00000000;
        12'b000000_000000: code<=32'b00000000_00000000_00000100_00000000;
        12'b000000_000010: code<=32'b00000000_00000000_00001000_00000000;
        12'b000000_000011: code<=32'b00000000_00000000_00010000_00000000;
        12'b000000_000100: code<=32'b00000000_00000000_00100000_00000000;
        12'b000000_000110: code<=32'b00000000_00000000_01000000_00000000;
        12'b000000_000111: code<=32'b00000000_00000000_10000000_00000000;
        12'b000000_001000: code<=32'b00000000_00000001_00000000_00000000;

        12'b001000_xxxxxx: code<=32'b00000000_00000010_00000000_00000000;
        12'b001001_xxxxxx: code<=32'b00000000_00000100_00000000_00000000;
        12'b001100_xxxxxx: code<=32'b00000000_00001000_00000000_00000000;
        12'b001101_xxxxxx: code<=32'b00000000_00010000_00000000_00000000;
        12'b001110_xxxxxx: code<=32'b00000000_00100000_00000000_00000000;
        12'b001111_xxxxxx: code<=32'b00000000_01000000_00000000_00000000;
        12'b100011_xxxxxx: code<=32'b00000000_10000000_00000000_00000000;
        12'b101011_xxxxxx: code<=32'b00000001_00000000_00000000_00000000;
        12'b000100_xxxxxx: code<=32'b00000010_00000000_00000000_00000000;
        12'b000101_xxxxxx: code<=32'b00000100_00000000_00000000_00000000;
        12'b001010_xxxxxx: code<=32'b00001000_00000000_00000000_00000000;
        12'b001011_xxxxxx: code<=32'b00010000_00000000_00000000_00000000;
        
        12'b000010_xxxxxx: code<=32'b00100000_00000000_00000000_00000000;
        12'b000011_xxxxxx: code<=32'b01000000_00000000_00000000_00000000;

        default: 
            code<=32'bz;
    endcase
end
    


endmodule //instrument_decoder